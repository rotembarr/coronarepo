////////////////////////////////////////////////////////////////////////////////
//
// File name    : mix_columns.sv
// Date Created : 13

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: The module to mix all the columns together.
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: 
//
////////////////////////////////////////////////////////////////////////////////

module mix_columns
(
	// Inputs and outputs

	input aes_model_pack::byte_table block_in,

	output aes_model_pack::byte_table mixed_block
);

	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	genvar i;

	// Generates a column mix for each column
	generate
		for (i = 0; i < aes_model_pack::COLUMN_COUNT; i++) begin : gen_columns
			mix_one_column moc_inst(
				.column      (block_in[i]),
				.mixed_column(mixed_block[i])
			);
		end
	endgenerate
endmodule // mix_columns