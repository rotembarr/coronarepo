// As the true top module contains QSYS files, and its problematic
// to simulate them, this tb is to simulate the top without the
// AES module. This testbench should be updated manually


module aes_top_tb ();



endmodule