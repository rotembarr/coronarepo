////////////////////////////////////////////////////////////////////////////////
//
// File name    : sub_bytes.sv
// Date Created : 14/8

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: Block sub bytes module
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: 
//
////////////////////////////////////////////////////////////////////////////////

module sub_bytes
(
	input aes_model_pack::byte_table plain_block,
	output aes_model_pack::byte_table sub_block
);
	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	always_comb begin : proc_sub
		for (int i = 0; i < aes_model_pack::COLUMN_COUNT; i++) begin
			for (int j = 0; j < aes_model_pack::COLUMN_SIZE_IN_BYTES; j++) begin
				
				// Transforms each byte to the one in the Sub bytes table
				sub_block[i][j] = aes_model_pack::SUB_BYTES_TABLE[plain_block[i][j]];	
			end
		end
	end
endmodule