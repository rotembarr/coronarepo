// single_port_ram.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module single_port_ram (
		input  wire         clk_clk,                        //                 clk.clk
		input  wire [5:0]   onchip_memory2_0_s1_address,    // onchip_memory2_0_s1.address
		input  wire         onchip_memory2_0_s1_clken,      //                    .clken
		input  wire         onchip_memory2_0_s1_chipselect, //                    .chipselect
		input  wire         onchip_memory2_0_s1_write,      //                    .write
		output wire [511:0] onchip_memory2_0_s1_readdata,   //                    .readdata
		input  wire [511:0] onchip_memory2_0_s1_writedata,  //                    .writedata
		input  wire [63:0]  onchip_memory2_0_s1_byteenable, //                    .byteenable
		input  wire [5:0]   onchip_memory2_0_s2_address,    // onchip_memory2_0_s2.address
		input  wire         onchip_memory2_0_s2_chipselect, //                    .chipselect
		input  wire         onchip_memory2_0_s2_clken,      //                    .clken
		input  wire         onchip_memory2_0_s2_write,      //                    .write
		output wire [511:0] onchip_memory2_0_s2_readdata,   //                    .readdata
		input  wire [511:0] onchip_memory2_0_s2_writedata,  //                    .writedata
		input  wire [63:0]  onchip_memory2_0_s2_byteenable, //                    .byteenable
		input  wire         reset_reset_n                   //               reset.reset_n
	);

	wire    rst_controller_reset_out_reset;     // rst_controller:reset_out -> onchip_memory2_0:reset
	wire    rst_controller_reset_out_reset_req; // rst_controller:reset_req -> onchip_memory2_0:reset_req

	single_port_ram_onchip_memory2_0 onchip_memory2_0 (
		.address     (onchip_memory2_0_s1_address),        //     s1.address
		.clken       (onchip_memory2_0_s1_clken),          //       .clken
		.chipselect  (onchip_memory2_0_s1_chipselect),     //       .chipselect
		.write       (onchip_memory2_0_s1_write),          //       .write
		.readdata    (onchip_memory2_0_s1_readdata),       //       .readdata
		.writedata   (onchip_memory2_0_s1_writedata),      //       .writedata
		.byteenable  (onchip_memory2_0_s1_byteenable),     //       .byteenable
		.address2    (onchip_memory2_0_s2_address),        //     s2.address
		.chipselect2 (onchip_memory2_0_s2_chipselect),     //       .chipselect
		.clken2      (onchip_memory2_0_s2_clken),          //       .clken
		.write2      (onchip_memory2_0_s2_write),          //       .write
		.readdata2   (onchip_memory2_0_s2_readdata),       //       .readdata
		.writedata2  (onchip_memory2_0_s2_writedata),      //       .writedata
		.byteenable2 (onchip_memory2_0_s2_byteenable),     //       .byteenable
		.clk         (clk_clk),                            //   clk1.clk
		.reset       (rst_controller_reset_out_reset),     // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
