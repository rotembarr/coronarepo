////////////////////////////////////////////////////////////////////////////////
//
// File name    : round_cipher_tb.sv
// Date Created : 14

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: Round cipher testbench
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: 
//
////////////////////////////////////////////////////////////////////////////////

module round_cipher_tb();
	///////////////////////////////////////////////////////////////////////////
	/////// Declarations //////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	logic clk = 1'b0;

	aes_model_pack::byte_table expected_output = {128'ha4686b029c9f5b6a7f35ea50f22b4349};

	aes_model_pack::byte_table state = {
		{8'h19, 8'ha0, 8'h9a, 8'he9},
		{8'h3d, 8'hf4, 8'hc6, 8'hf8},
		{8'he3, 8'he2, 8'h8d, 8'h48},
		{8'hbe, 8'h2b, 8'h2a, 8'h08}
	};
	aes_model_pack::byte_table round_key = {
		{8'ha0, 8'h88, 8'h23, 8'h2a},
		{8'hfa, 8'h54, 8'ha3, 8'h6c},
		{8'hfe, 8'h2c, 8'h39, 8'h76},
		{8'h17, 8'hb1, 8'h39, 8'h05}
	};

	aes_model_pack::byte_table cipher_block;

	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	always
	begin
		#aes_const_pack::CLK_FREQ clk =~clk;
	end

	initial	begin
		#20ns;
		@(posedge clk);
		$display("%h",cipher_block);
		assert (expected_output == cipher_block) begin
			$display("Correct output");
		end
		else begin
			$display("Wrong");
		end
		$finish();
	end

	///////////////////////////////////////////////////////////////////////////
	/////// Instantiations ////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	round_cipher dut(
		.state       (state),
		.round_key   (round_key),
		.last_round  (1'b0),
		.cipher_state(cipher_block)
	);
	
endmodule // round_cipher_tb