////////////////////////////////////////////////////////////////////////////////
//
// File name    : sub_bytes_tb.sv
// Date Created : 14

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: Sub bytes testbench
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: 
//
////////////////////////////////////////////////////////////////////////////////

module sub_bytes_tb();
	///////////////////////////////////////////////////////////////////////////
	/////// Declarations //////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	logic clk = 1'b0;

	aes_model_pack::byte_table pre_sub = {
		{8'h19, 8'ha0, 8'h9a, 8'he9},
		{8'h3d, 8'hf4, 8'hc6, 8'hf8},
		{8'he3, 8'he2, 8'h8d, 8'h48},
		{8'hbe, 8'h2b, 8'h2a, 8'h08}
	};

	aes_model_pack::byte_table post_sub;

	aes_model_pack::byte_table result = 128'hd4e0b81e27bfb44111985d52aef1e530;


	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	sub_bytes dut(
		.plain_block(pre_sub),
		.sub_block  (post_sub)
	);

	always begin
		#aes_const_pack::CLK_FREQ clk = ~clk;
	end

	initial begin
		#20ns;
		@(posedge clk);
		$display("%h",pre_sub);
		$display("%h",post_sub);
		assert (post_sub == result);
		$finish();
	end

endmodule