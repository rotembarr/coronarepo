////////////////////////////////////////////////////////////////////////////////
//
// File name    : shift_rows_tb.sv
// Date Created : 14

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: Testbench for shift rows
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: 
//
////////////////////////////////////////////////////////////////////////////////

module shift_rows_tb();
	///////////////////////////////////////////////////////////////////////////
	/////// Declarations //////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	logic clk = 1'b0;

	aes_model_pack::byte_table pre_shift = {
		{8'h15,	8'h14,	8'h13,	8'h12	},
		{8'h11,	8'h10,	8'h9,	8'h8	},
		{8'h7,	8'h6,	8'h5,	8'h4 	},
		{8'h3,	8'h2,	8'h1,	8'h0 	}
	};

	aes_model_pack::byte_table after_shift;

	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	
	always begin
		#aes_const_pack::CLK_FREQ clk = ~clk;
	end

	initial begin
		#20ns;
		@(posedge clk);
		$display("%h", pre_shift);
		$display("%h", after_shift);
		$finish();
	end

	///////////////////////////////////////////////////////////////////////////
	/////// Instantiations ////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	shift_rows dut(
		.state      (pre_shift),
		.shift_block(after_shift)
	);

endmodule