///////////////////////////////////////////////
// This module's purpose is to allow future  //
// debug access using the registers. 		 //
///////////////////////////////////////////////

module registers_controller 
#(
	parameter int COUNTER_SIZE = 32
)
(
	// General
	input logic clk,
	input logic rst_n,
	
	// Avalon-mm
);

endmodule