////////////////////////////////////////////////////////////////////////////////
//
// File name    : key_warm_tb.sv
// Date Created : 21

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: Key warm testbench
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: 
//
////////////////////////////////////////////////////////////////////////////////

module key_warm_tb();
	///////////////////////////////////////////////////////////////////////////
	/////// Declarations //////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	logic clk = 1'b0;
	logic rst = 1'b0;

	// Key input
	aes_model_pack::byte_table key = { 128'h2b7e151628aed2a6abf7158809cf4f3c };
	//aes_model_pack::byte_table key = '0;

	// Key signals
	logic warm_key  = 1'b0;
	logic reset_key = 1'b0;

	// Key output
	aes_model_pack::byte_table key_round;
	aes_model_pack::byte_table expected_output = { 128'hd014f9a8c9ee2589e13f0cc8b6630ca6 };


	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	always begin
		#aes_model_pack::CLK_FREQ clk = ~clk;
	end

	initial begin

		// Reset process
		#20ns;
		@(posedge clk);
		rst = 1'b1;

		// Start key warm
		@(posedge clk);
		warm_key = 1'b1;

		// Key process
		repeat (aes_model_pack::ROUND_COUNT) begin
			@(posedge clk);
		end

		warm_key = 1'b0;

		@(posedge clk);
		assert (key_round == expected_output) begin
			$display("ok");
		end else begin
			$display("not ok");
			$display("got %p", key_round);
		end
		$finish();
	end

	///////////////////////////////////////////////////////////////////////////
	/////// Instantiations ////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	key_warm dut (
		.clk(clk),
		.rst(rst),
		.key(key),
		.warm_key (warm_key ),
		.key_round(key_round)
	);

endmodule