////////////////////////////////////////////////////////////////////////////////
//
// File name    : mix_one_column_tb.sv
// Date Created : 14

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: Testbench for mix_one_column
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: Using inputs that their output is known to check if the calculation
//			 is correct.
//
////////////////////////////////////////////////////////////////////////////////

module mix_one_column_tb();
	///////////////////////////////////////////////////////////////////////////
	/////// Localparams ///////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	localparam int INPUT_COLUMNS = 4;

	///////////////////////////////////////////////////////////////////////////
	/////// Declarations //////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	logic clk 	  																	= 1'b0;
	logic [aes_model_pack::COLUMN_SIZE_IN_BYTES-1:0][$bits(byte)-1:0] input_column;
	logic [aes_model_pack::COLUMN_SIZE_IN_BYTES-1:0][$bits(byte)-1:0] output_column;
	int  															  index 		= 0;

	//Selected inputs for the columns, as the output is known
	logic [INPUT_COLUMNS-1:0][aes_model_pack::COLUMN_SIZE_IN_BYTES-1:0][$bits(byte)-1:0] columns = {
		{8'hf2, 8'h0a, 8'h22, 8'h5c}, //Should output [9f,dc,58,9d]
		{8'hdb, 8'he0, 8'hb8, 8'h1e}, //Should output [8e,4d,a1,bc]
		{8'h01, 8'h01, 8'h01, 8'h01}, //Should output the same
		{8'hd4, 8'hd4, 8'hd4, 8'hd5}  //Should output [d5,d5,d7,d6]
	};


	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	always
    begin
        #test_pack::CLK_FREQ clk = ~clk;
    end


	initial	begin
		index = 0;
		input_column <= columns[index];
		#20ns;
		repeat (INPUT_COLUMNS + 1) begin
			index <= index + 1;
			$display("input %h", input_column);
			$display("output %h", output_column);
			@(posedge clk);
			input_column <= columns[index];
		end
		$finish();
	end

	///////////////////////////////////////////////////////////////////////////
	/////// Instantiations ////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	mix_one_column dut_inst(
		.column      (input_column),
		.mixed_column(output_column)
	);
endmodule // mix_one_column_tb