////////////////////////////////////////////////////////////////////////////////
//
// File name    : round_cipher.sv
// Date Created : 14

//
////////////////////////////////////////////////////////////////////////////////
//
// Description: The module for the round process
//
////////////////////////////////////////////////////////////////////////////////
//
// Comments: 
//
////////////////////////////////////////////////////////////////////////////////

module round_cipher
(
	// Inputs and outputs

	input aes_model_pack::byte_table state,
	input aes_model_pack::byte_table round_key,
	input logic  	  				 last_round,

	output aes_model_pack::byte_table cipher_state
);
	///////////////////////////////////////////////////////////////////////////
	/////// Declarations //////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	aes_model_pack::byte_table sub_block, shift_block, mixed_block, sel_block;

	///////////////////////////////////////////////////////////////////////////
	/////// Logic /////////////////////////////////////////////////////////////
	///////////////////////////////////////////////////////////////////////////

	sub_bytes sub_bytes_inst(
		.plain_block(state), // Input
		.sub_block  (sub_block) // Output
	);

	shift_rows shift_rows_inst(
		.state      (sub_block), // Input
		.shift_block(shift_block) // Output
	);

	mix_columns mix_columns_inst(
		.block_in   (shift_block), // Input
		.mixed_block(mixed_block) // Output
	);

	assign sel_block = (last_round) ? shift_block : mixed_block;
	assign cipher_state = sel_block ^ round_key;

endmodule // round_cipher